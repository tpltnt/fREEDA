Simple RC network

r1 1 2 500
c1 0 2 5p 
* c1 0 2 5p ic=2V
vin 1 0 pulse (0 1.5 4ns 3ns 5ns 2ns 17ns)
.tran 500ps 34ns 
*.dc vin 0 0.1 0.001 
*.print dc v(1) v(2)
* .options numdgt=7
.Four 58.8235MegHz V(1) V(2)
.print tran v(1) v(2) i(vin)
.end
