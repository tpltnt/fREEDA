RLC filter
*
* `Short' input so that it does not form
* part of the output impedance
*Vin 1 0 AC 0V
Vin 1 0 AC 1V
*
R1 1 2 15Ohm
L1 2 3 50mH
C1 3 0 1.5uF
*
* AC statement just defines frequency range
.AC dec 20 100Hz 10kHz
*
* Noise analysis at Node 3 with respect of Vin
.noise V(3) Vin 10
*
* Measure output impedance with a current source
* Iout 0 3 AC 1
*
* Measure Zout:
*.print AC VM(3)
*
*
.print NOISE INOISE

.end
